
module kernel (
	clk_clk,
	pio_nco_phi_export,
	reset_reset_n);	

	input		clk_clk;
	output	[31:0]	pio_nco_phi_export;
	input		reset_reset_n;
endmodule
